   // RANDOM GENERATOR of A and B
class RCSG;

	rand bit [sys_iff.A_bits -1:0]  A_;
    rand bit [sys_iff.B_bits -1:0]  B_;

endclass