   // RANDOM GENERATOR of A and B
    
    class RCSG;

        system_iff sys_iff;

	    rand bit [sys_iff.A_bits -1:0]  sys_iff.A;
        rand bit [sys_iff.B_bits -1:0]  sys_iff.B;


    endclass