`include "memory.sv"
`include "register_bank.sv"

/**
    @brief Top level entity for the RISC-V processor
*/
module top_processor(

);

// Instanciate the data path

// Instanciate the control module





endmodule
