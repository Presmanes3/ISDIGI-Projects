class scoreboard;

system_iff sys_iff;


task multiply(reg A,reg B);
    
endtask

task compare_outputs(reg ideal_result, reg real_result);

endtask
endclass