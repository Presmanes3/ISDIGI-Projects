module alu_controller(

    input   []      alu_option;  
    output  [3:0]   alu_operation;
);




endmodule