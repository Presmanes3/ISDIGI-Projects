
module sum_shift_based_multiplier (
    
);


    
endmodule