module clear_pipeline_designator (
    segmented_interface wires
);


    
endmodule