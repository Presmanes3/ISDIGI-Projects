`include "memory.sv"
`include "register_bank.sv"

/**
    @brief Top level entity for the RISC-V processor
*/
module core(

);

// Instanciate the data path

// Instanciate the control module





endmodule
