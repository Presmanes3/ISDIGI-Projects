module main_controller(

    
);





endmodule