module hazard_detection_unit_designator (
    segmented_interface wires
);
    
endmodule