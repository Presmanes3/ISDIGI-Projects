   // RANDOM GENERATOR of A and B
class RCSG;

	rand bit [testbench.sys_iff.A_bits -1:0]  A_;
    rand bit [testbench.sys_iff.B_bits -1:0]  B_;

endclass