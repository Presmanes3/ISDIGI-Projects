class scoreboard;

system_iff sys_iff;


task multiply();
    
endtask

task compare_outputs();

endtask

endclass