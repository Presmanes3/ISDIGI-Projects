module data_forwarding_designator (
    segmented_interface wires
);


    
endmodule