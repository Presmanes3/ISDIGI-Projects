module testbench(
    
);
    

    
endmodule